----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.all;

use IEEE.NUMERIC_STD.all;
use IEEE.MATH_REAL.all;                 -- for simulation

entity tb_math is
--  Port ( );
end tb_math;

architecture Behavioral of tb_math is
  signal clk             : std_logic                     := '0';
  signal reset           : std_logic                     := '0';
  signal start           : std_logic                     := '0';
  signal done            : std_logic                     := '0';
  signal a               : std_logic_vector(39 downto 0) := (others => '0');
  signal b               : std_logic_vector(39 downto 0) := (others => '0');
  signal c               : std_logic_vector(39 downto 0) := (others => '0');
  signal op              : std_logic_vector(3 downto 0) := (others => '0');
  signal err             : std_logic                     := '0';
  signal simulation_done : boolean                       := false;
begin

  r1 : entity work.kmath(Behavioral) port map
    (
      i_clk       => clk,
      i_reset     => reset,
      i_start     => start,
      i_a         => a,
      i_b         => b,
      i_op        => op,
      o_done      => done,
      o_c         => c,
      o_err       => err
      );

  clk <= not clk after 5 ns when not simulation_done else '0';

  p : process is
    variable per       : integer := 100;
    variable failures  : integer := 0;
    variable err_count : integer := 0;
    variable vec_fails : integer := 0;
    variable runs      : integer := 0;

    -- note: due to restriciton in vhdl ints we can't actually check the
    -- values from 2**31 to 2**32-1 we just assume they work
    procedure run(iop : std_logic_vector(3 downto 0);
                  aa, bb : std_logic_vector(39 downto 0)) is
      variable expected : real;
      variable result   : real;
      variable realp    : real;
    begin
      wait until rising_edge(clk);
      op(3 downto 0) <= iop;
      a(39 downto 0) <= aa;
      b(39 downto 0) <= bb;
      wait until rising_edge(clk);
      start          <= '1';
      wait until rising_edge(clk);
      start          <= '0';
      if done = '0' then
        wait until rising_edge(clk);
      end if;

      wait until done = '1';
      wait until rising_edge(clk);

      if err = '1' then
        err_count := err_count + 1;
        report "DUT err reported" severity warning;
      end if;


      runs := runs + 1;

    end;

    procedure run_uint(iop : std_logic_vector(3 downto 0);
                       aa, bb : integer range 0 to 2**31 - 1) is
    begin
      run( iop => iop,
           aa => std_logic_vector(to_unsigned(aa, 40)),
           bb => std_logic_vector(to_unsigned(bb, 40)));
    end;

    -- run and expect output cc
    procedure kvec(iop : std_logic_vector(3 downto 0);
                       aa, bb, cc : std_logic_vector(39 downto 0)) is
    begin
      run( iop => iop,aa => aa, bb => bb);

      if c /= cc then
        vec_fails := vec_fails + 1;
        report "DUT vector fail reported" severity failure;
      end if;
    end;

    

  begin
    wait for 5 ns;

    wait until rising_edge(clk);
    reset <= '1';
    wait until rising_edge(clk);
    reset <= '0';

    run( "0000", x"ff_ffff_fff6", x"00_0000_0000");

    run( "0001",               c, x"00_0000_0000");
    
    
    run_uint( "0000", 666, 22);                   -- 0x029a, 0x0016
    run_uint( "0000", 666, 22);                   -- 0x029a, 0x0016

    -- test out expected problematic inputs: 0,1,2,3 and very large values
    -- we expect at least some of these to trigger the range error
    err_count := 0;
    run_uint( "0000", 0, 0);
    run_uint( "0000", 1, 0);
    run_uint( "0000", 256, 0);

    -- the "C" code produces a KVEC procedure call each time the unit
    -- is called, so we can just cut and paste all these in using (from bash)
    -- for P in tc/*txt; do grep -h KVEC $P ; done

KVEC(x"4",x"40d0000000", x"40d0000000", x"4150000000");
KVEC(x"4",x"0000000000", x"7fffffffff", x"7fffffffff");
KVEC(x"2",x"7fffffffff", x"7fffffffff", x"7fffffffff");
KVEC(x"0",x"fffffffff6", x"0000000000", x"c150000000");
KVEC(x"1",x"c150000000", x"0000000000", x"fffffffff6");
KVEC(x"0",x"fffffffff7", x"0000000000", x"c148000000");
KVEC(x"1",x"c148000000", x"0000000000", x"fffffffff7");
KVEC(x"0",x"fffffffff8", x"0000000000", x"c140000000");
KVEC(x"1",x"c140000000", x"0000000000", x"fffffffff8");
KVEC(x"0",x"fffffffff9", x"0000000000", x"c0f0000000");
KVEC(x"1",x"c0f0000000", x"0000000000", x"fffffffff9");
KVEC(x"4",x"7f80000000", x"40d0000000", x"7f80000000");
KVEC(x"0",x"fffffffffa", x"0000000000", x"c0e0000000");
KVEC(x"1",x"c0e0000000", x"0000000000", x"fffffffffa");
KVEC(x"0",x"fffffffffb", x"0000000000", x"c0d0000000");
KVEC(x"1",x"c0d0000000", x"0000000000", x"fffffffffb");
KVEC(x"0",x"fffffffffc", x"0000000000", x"c0c0000000");
KVEC(x"1",x"c0c0000000", x"0000000000", x"fffffffffc");
KVEC(x"0",x"fffffffffd", x"0000000000", x"c060000000");
KVEC(x"1",x"c060000000", x"0000000000", x"fffffffffd");
KVEC(x"0",x"fffffffffe", x"0000000000", x"c040000000");
KVEC(x"1",x"c040000000", x"0000000000", x"fffffffffe");
KVEC(x"4",x"7f80000000", x"0000000000", x"7f80000000");
KVEC(x"0",x"ffffffffff", x"0000000000", x"bfc0000000");
KVEC(x"1",x"bfc0000000", x"0000000000", x"ffffffffff");
KVEC(x"0",x"0000000000", x"0000000000", x"0000000000");
KVEC(x"1",x"0000000000", x"0000000000", x"0000000000");
KVEC(x"0",x"0000000001", x"0000000000", x"3fc0000000");
KVEC(x"1",x"3fc0000000", x"0000000000", x"0000000001");
KVEC(x"0",x"0000000002", x"0000000000", x"4040000000");
KVEC(x"1",x"4040000000", x"0000000000", x"0000000002");
KVEC(x"0",x"0000000003", x"0000000000", x"4060000000");
KVEC(x"1",x"4060000000", x"0000000000", x"0000000003");
KVEC(x"4",x"7f80000000", x"7f80000000", x"7f80000000");
KVEC(x"0",x"0000000004", x"0000000000", x"40c0000000");
KVEC(x"1",x"40c0000000", x"0000000000", x"0000000004");
KVEC(x"0",x"0000000005", x"0000000000", x"40d0000000");
KVEC(x"1",x"40d0000000", x"0000000000", x"0000000005");
KVEC(x"0",x"0000000006", x"0000000000", x"40e0000000");
KVEC(x"1",x"40e0000000", x"0000000000", x"0000000006");
KVEC(x"0",x"0000000007", x"0000000000", x"40f0000000");
KVEC(x"1",x"40f0000000", x"0000000000", x"0000000007");
KVEC(x"0",x"0000000008", x"0000000000", x"4140000000");
KVEC(x"1",x"4140000000", x"0000000000", x"0000000008");
KVEC(x"4",x"7f80000000", x"ff80000000", x"7fffffffff");
KVEC(x"0",x"0000000009", x"0000000000", x"4148000000");
KVEC(x"1",x"4148000000", x"0000000000", x"0000000009");
KVEC(x"0",x"0000000002", x"0000000000", x"4040000000");
KVEC(x"1",x"4040000000", x"0000000000", x"0000000002");
KVEC(x"0",x"0000000004", x"0000000000", x"40c0000000");
KVEC(x"1",x"40c0000000", x"0000000000", x"0000000004");
KVEC(x"0",x"0000000008", x"0000000000", x"4140000000");
KVEC(x"1",x"4140000000", x"0000000000", x"0000000008");
KVEC(x"0",x"0000000010", x"0000000000", x"41c0000000");
KVEC(x"1",x"41c0000000", x"0000000000", x"0000000010");
KVEC(x"4",x"7f80000000", x"7fffffffff", x"7fffffffff");
KVEC(x"0",x"0000000020", x"0000000000", x"4240000000");
KVEC(x"1",x"4240000000", x"0000000000", x"0000000020");
KVEC(x"0",x"0000000040", x"0000000000", x"42c0000000");
KVEC(x"1",x"42c0000000", x"0000000000", x"0000000040");
KVEC(x"0",x"0000000080", x"0000000000", x"4340000000");
KVEC(x"1",x"4340000000", x"0000000000", x"0000000080");
KVEC(x"0",x"0000000100", x"0000000000", x"43c0000000");
KVEC(x"1",x"43c0000000", x"0000000000", x"0000000100");
KVEC(x"0",x"0000000200", x"0000000000", x"4440000000");
KVEC(x"1",x"4440000000", x"0000000000", x"0000000200");
KVEC(x"4",x"ff80000000", x"40d0000000", x"ff80000000");
KVEC(x"0",x"0000000400", x"0000000000", x"44c0000000");
KVEC(x"1",x"44c0000000", x"0000000000", x"0000000400");
KVEC(x"0",x"0000000800", x"0000000000", x"4540000000");
KVEC(x"1",x"4540000000", x"0000000000", x"0000000800");
KVEC(x"0",x"0000001000", x"0000000000", x"45c0000000");
KVEC(x"1",x"45c0000000", x"0000000000", x"0000001000");
KVEC(x"0",x"0000002000", x"0000000000", x"4640000000");
KVEC(x"1",x"4640000000", x"0000000000", x"0000002000");
KVEC(x"0",x"0000004000", x"0000000000", x"46c0000000");
KVEC(x"1",x"46c0000000", x"0000000000", x"0000004000");
KVEC(x"4",x"ff80000000", x"0000000000", x"ff80000000");
KVEC(x"0",x"0000008000", x"0000000000", x"4740000000");
KVEC(x"1",x"4740000000", x"0000000000", x"0000008000");
KVEC(x"0",x"0000010000", x"0000000000", x"47c0000000");
KVEC(x"1",x"47c0000000", x"0000000000", x"0000010000");
KVEC(x"0",x"0000020000", x"0000000000", x"4840000000");
KVEC(x"1",x"4840000000", x"0000000000", x"0000020000");
KVEC(x"0",x"0000040000", x"0000000000", x"48c0000000");
KVEC(x"1",x"48c0000000", x"0000000000", x"0000040000");
KVEC(x"0",x"0000080000", x"0000000000", x"4940000000");
KVEC(x"1",x"4940000000", x"0000000000", x"0000080000");
KVEC(x"4",x"ff80000000", x"7f80000000", x"7fffffffff");
KVEC(x"0",x"0000100000", x"0000000000", x"49c0000000");
KVEC(x"1",x"49c0000000", x"0000000000", x"0000100000");
KVEC(x"0",x"0000200000", x"0000000000", x"4a40000000");
KVEC(x"1",x"4a40000000", x"0000000000", x"0000200000");
KVEC(x"0",x"0000400000", x"0000000000", x"4ac0000000");
KVEC(x"1",x"4ac0000000", x"0000000000", x"0000400000");
KVEC(x"0",x"0000800000", x"0000000000", x"4b40000000");
KVEC(x"1",x"4b40000000", x"0000000000", x"0000800000");
KVEC(x"0",x"0001000000", x"0000000000", x"4bc0000000");
KVEC(x"1",x"4bc0000000", x"0000000000", x"0001000000");
KVEC(x"4",x"ff80000000", x"ff80000000", x"ff80000000");
KVEC(x"0",x"0002000000", x"0000000000", x"4c40000000");
KVEC(x"1",x"4c40000000", x"0000000000", x"0002000000");
KVEC(x"0",x"0004000000", x"0000000000", x"4cc0000000");
KVEC(x"1",x"4cc0000000", x"0000000000", x"0004000000");
KVEC(x"0",x"0008000000", x"0000000000", x"4d40000000");
KVEC(x"1",x"4d40000000", x"0000000000", x"0008000000");
KVEC(x"0",x"0010000000", x"0000000000", x"4dc0000000");
KVEC(x"1",x"4dc0000000", x"0000000000", x"0010000000");
KVEC(x"0",x"0020000000", x"0000000000", x"4e40000000");
KVEC(x"1",x"4e40000000", x"0000000000", x"0020000000");
KVEC(x"4",x"40d0000000", x"0000000000", x"40d0000000");
KVEC(x"4",x"ff80000000", x"7fffffffff", x"7fffffffff");
KVEC(x"0",x"0040000000", x"0000000000", x"4ec0000000");
KVEC(x"1",x"4ec0000000", x"0000000000", x"0040000000");
KVEC(x"1",x"c040000000", x"0000000000", x"fffffffffe");
KVEC(x"0",x"fffffffffe", x"0000000000", x"c040000000");
KVEC(x"1",x"c0c0000000", x"0000000000", x"fffffffffc");
KVEC(x"0",x"fffffffffc", x"0000000000", x"c0c0000000");
KVEC(x"1",x"c140000000", x"0000000000", x"fffffffff8");
KVEC(x"0",x"fffffffff8", x"0000000000", x"c140000000");
KVEC(x"1",x"c1c0000000", x"0000000000", x"fffffffff0");
KVEC(x"0",x"fffffffff0", x"0000000000", x"c1c0000000");
KVEC(x"4",x"7fffffffff", x"40d0000000", x"7fffffffff");
KVEC(x"1",x"c240000000", x"0000000000", x"ffffffffe0");
KVEC(x"0",x"ffffffffe0", x"0000000000", x"c240000000");
KVEC(x"1",x"c2c0000000", x"0000000000", x"ffffffffc0");
KVEC(x"0",x"ffffffffc0", x"0000000000", x"c2c0000000");
KVEC(x"1",x"c340000000", x"0000000000", x"ffffffff80");
KVEC(x"0",x"ffffffff80", x"0000000000", x"c340000000");
KVEC(x"1",x"c3c0000000", x"0000000000", x"ffffffff00");
KVEC(x"0",x"ffffffff00", x"0000000000", x"c3c0000000");
KVEC(x"1",x"c440000000", x"0000000000", x"fffffffe00");
KVEC(x"0",x"fffffffe00", x"0000000000", x"c440000000");
KVEC(x"4",x"7fffffffff", x"0000000000", x"7fffffffff");
KVEC(x"1",x"c4c0000000", x"0000000000", x"fffffffc00");
KVEC(x"0",x"fffffffc00", x"0000000000", x"c4c0000000");
KVEC(x"1",x"c540000000", x"0000000000", x"fffffff800");
KVEC(x"0",x"fffffff800", x"0000000000", x"c540000000");
KVEC(x"1",x"c5c0000000", x"0000000000", x"fffffff000");
KVEC(x"0",x"fffffff000", x"0000000000", x"c5c0000000");
KVEC(x"1",x"c640000000", x"0000000000", x"ffffffe000");
KVEC(x"0",x"ffffffe000", x"0000000000", x"c640000000");
KVEC(x"1",x"c6c0000000", x"0000000000", x"ffffffc000");
KVEC(x"0",x"ffffffc000", x"0000000000", x"c6c0000000");
KVEC(x"4",x"7fffffffff", x"7f80000000", x"7fffffffff");
KVEC(x"1",x"c740000000", x"0000000000", x"ffffff8000");
KVEC(x"0",x"ffffff8000", x"0000000000", x"c740000000");
KVEC(x"1",x"c7c0000000", x"0000000000", x"ffffff0000");
KVEC(x"0",x"ffffff0000", x"0000000000", x"c7c0000000");
KVEC(x"1",x"c840000000", x"0000000000", x"fffffe0000");
KVEC(x"0",x"fffffe0000", x"0000000000", x"c840000000");
KVEC(x"1",x"c8c0000000", x"0000000000", x"fffffc0000");
KVEC(x"0",x"fffffc0000", x"0000000000", x"c8c0000000");
KVEC(x"1",x"c940000000", x"0000000000", x"fffff80000");
KVEC(x"0",x"fffff80000", x"0000000000", x"c940000000");
KVEC(x"4",x"7fffffffff", x"ff80000000", x"7fffffffff");
KVEC(x"1",x"c9c0000000", x"0000000000", x"fffff00000");
KVEC(x"0",x"fffff00000", x"0000000000", x"c9c0000000");
KVEC(x"1",x"ca40000000", x"0000000000", x"ffffe00000");
KVEC(x"0",x"ffffe00000", x"0000000000", x"ca40000000");
KVEC(x"1",x"cac0000000", x"0000000000", x"ffffc00000");
KVEC(x"0",x"ffffc00000", x"0000000000", x"cac0000000");
KVEC(x"1",x"cb40000000", x"0000000000", x"ffff800000");
KVEC(x"0",x"ffff800000", x"0000000000", x"cb40000000");
KVEC(x"1",x"cbc0000000", x"0000000000", x"ffff000000");
KVEC(x"0",x"ffff000000", x"0000000000", x"cbc0000000");
KVEC(x"4",x"7fffffffff", x"7fffffffff", x"7fffffffff");
KVEC(x"1",x"cc40000000", x"0000000000", x"fffe000000");
KVEC(x"0",x"fffe000000", x"0000000000", x"cc40000000");
KVEC(x"1",x"ccc0000000", x"0000000000", x"fffc000000");
KVEC(x"0",x"fffc000000", x"0000000000", x"ccc0000000");
KVEC(x"1",x"cd40000000", x"0000000000", x"fff8000000");
KVEC(x"0",x"fff8000000", x"0000000000", x"cd40000000");
KVEC(x"1",x"cdc0000000", x"0000000000", x"fff0000000");
KVEC(x"0",x"fff0000000", x"0000000000", x"cdc0000000");
KVEC(x"1",x"ce40000000", x"0000000000", x"ffe0000000");
KVEC(x"0",x"ffe0000000", x"0000000000", x"ce40000000");
KVEC(x"5",x"40d0000000", x"40d0000000", x"0000000000");
KVEC(x"1",x"cec0000000", x"0000000000", x"ffc0000000");
KVEC(x"0",x"ffc0000000", x"0000000000", x"cec0000000");
KVEC(x"1",x"cf40000000", x"0000000000", x"ff80000000");
KVEC(x"0",x"ff80000000", x"0000000000", x"cf40000000");
KVEC(x"2",x"0000000000", x"4168000000", x"0000000000");
KVEC(x"2",x"447bc00000", x"0000000000", x"7f80000000");
KVEC(x"2",x"42e4000000", x"4168000000", x"40fb13b13a");
KVEC(x"2",x"c150000000", x"c150000000", x"3fc0000000");
KVEC(x"2",x"c150000000", x"c148000000", x"3fc71c71c7");
KVEC(x"2",x"c150000000", x"c140000000", x"3fd0000000");
KVEC(x"5",x"40d0000000", x"0000000000", x"40d0000000");
KVEC(x"2",x"c150000000", x"c0f0000000", x"3fdb6db6da");
KVEC(x"2",x"c150000000", x"c0e0000000", x"3feaaaaaaa");
KVEC(x"2",x"c150000000", x"c0d0000000", x"4040000000");
KVEC(x"2",x"c150000000", x"c0c0000000", x"4050000000");
KVEC(x"2",x"c150000000", x"c060000000", x"406aaaaaaa");
KVEC(x"2",x"c150000000", x"c040000000", x"40d0000000");
KVEC(x"2",x"c150000000", x"bfc0000000", x"4150000000");
KVEC(x"2",x"c150000000", x"0000000000", x"ff80000000");
KVEC(x"2",x"c150000000", x"3fc0000000", x"c150000000");
KVEC(x"2",x"c150000000", x"4040000000", x"c0d0000000");
KVEC(x"5",x"40d0000000", x"7f80000000", x"ff80000000");
KVEC(x"2",x"c150000000", x"4060000000", x"c06aaaaaaa");
KVEC(x"2",x"c150000000", x"40c0000000", x"c050000000");
KVEC(x"2",x"c150000000", x"40d0000000", x"c040000000");
KVEC(x"2",x"c150000000", x"40e0000000", x"bfeaaaaaaa");
KVEC(x"2",x"c150000000", x"40f0000000", x"bfdb6db6da");
KVEC(x"2",x"c150000000", x"4140000000", x"bfd0000000");
KVEC(x"2",x"c150000000", x"4148000000", x"bfc71c71c7");
KVEC(x"2",x"c148000000", x"c150000000", x"3f73333332");
KVEC(x"2",x"c148000000", x"c148000000", x"3fc0000000");
KVEC(x"2",x"c148000000", x"c140000000", x"3fc8000000");
KVEC(x"5",x"40d0000000", x"ff80000000", x"7f80000000");
KVEC(x"2",x"c148000000", x"c0f0000000", x"3fd2492492");
KVEC(x"2",x"c148000000", x"c0e0000000", x"3fe0000000");
KVEC(x"2",x"c148000000", x"c0d0000000", x"3ff3333332");
KVEC(x"2",x"c148000000", x"c0c0000000", x"4048000000");
KVEC(x"2",x"c148000000", x"c060000000", x"4060000000");
KVEC(x"2",x"c148000000", x"c040000000", x"40c8000000");
KVEC(x"2",x"c148000000", x"bfc0000000", x"4148000000");
KVEC(x"2",x"c148000000", x"0000000000", x"ff80000000");
KVEC(x"2",x"c148000000", x"3fc0000000", x"c148000000");
KVEC(x"2",x"c148000000", x"4040000000", x"c0c8000000");
KVEC(x"4",x"40d0000000", x"7f80000000", x"7f80000000");
KVEC(x"5",x"40d0000000", x"7fffffffff", x"7fffffffff");
KVEC(x"2",x"c148000000", x"4060000000", x"c060000000");
KVEC(x"2",x"c148000000", x"40c0000000", x"c048000000");
KVEC(x"2",x"c148000000", x"40d0000000", x"bff3333332");
KVEC(x"2",x"c148000000", x"40e0000000", x"bfe0000000");
KVEC(x"2",x"c148000000", x"40f0000000", x"bfd2492492");
KVEC(x"2",x"c148000000", x"4140000000", x"bfc8000000");
KVEC(x"2",x"c148000000", x"4148000000", x"bfc0000000");
KVEC(x"2",x"c140000000", x"c150000000", x"3f66666666");
KVEC(x"2",x"c140000000", x"c148000000", x"3f71c71c70");
KVEC(x"2",x"c140000000", x"c140000000", x"3fc0000000");
KVEC(x"5",x"0000000000", x"40d0000000", x"c0d0000000");
KVEC(x"2",x"c140000000", x"c0f0000000", x"3fc9249248");
KVEC(x"2",x"c140000000", x"c0e0000000", x"3fd5555554");
KVEC(x"2",x"c140000000", x"c0d0000000", x"3fe6666666");
KVEC(x"2",x"c140000000", x"c0c0000000", x"4040000000");
KVEC(x"2",x"c140000000", x"c060000000", x"4055555554");
KVEC(x"2",x"c140000000", x"c040000000", x"40c0000000");
KVEC(x"2",x"c140000000", x"bfc0000000", x"4140000000");
KVEC(x"2",x"c140000000", x"0000000000", x"ff80000000");
KVEC(x"2",x"c140000000", x"3fc0000000", x"c140000000");
KVEC(x"2",x"c140000000", x"4040000000", x"c0c0000000");
KVEC(x"5",x"0000000000", x"0000000000", x"0000000000");
KVEC(x"2",x"c140000000", x"4060000000", x"c055555554");
KVEC(x"2",x"c140000000", x"40c0000000", x"c040000000");
KVEC(x"2",x"c140000000", x"40d0000000", x"bfe6666666");
KVEC(x"2",x"c140000000", x"40e0000000", x"bfd5555554");
KVEC(x"2",x"c140000000", x"40f0000000", x"bfc9249248");
KVEC(x"2",x"c140000000", x"4140000000", x"bfc0000000");
KVEC(x"2",x"c140000000", x"4148000000", x"bf71c71c70");
KVEC(x"2",x"c0f0000000", x"c150000000", x"3f59999999");
KVEC(x"2",x"c0f0000000", x"c148000000", x"3f638e38e3");
KVEC(x"2",x"c0f0000000", x"c140000000", x"3f70000000");
KVEC(x"5",x"0000000000", x"7f80000000", x"ff80000000");
KVEC(x"2",x"c0f0000000", x"c0f0000000", x"3fc0000000");
KVEC(x"2",x"c0f0000000", x"c0e0000000", x"3fcaaaaaaa");
KVEC(x"2",x"c0f0000000", x"c0d0000000", x"3fd9999999");
KVEC(x"2",x"c0f0000000", x"c0c0000000", x"3ff0000000");
KVEC(x"2",x"c0f0000000", x"c060000000", x"404aaaaaaa");
KVEC(x"2",x"c0f0000000", x"c040000000", x"4070000000");
KVEC(x"2",x"c0f0000000", x"bfc0000000", x"40f0000000");
KVEC(x"2",x"c0f0000000", x"0000000000", x"ff80000000");
KVEC(x"2",x"c0f0000000", x"3fc0000000", x"c0f0000000");
KVEC(x"2",x"c0f0000000", x"4040000000", x"c070000000");
KVEC(x"5",x"0000000000", x"ff80000000", x"7f80000000");
KVEC(x"2",x"c0f0000000", x"4060000000", x"c04aaaaaaa");
KVEC(x"2",x"c0f0000000", x"40c0000000", x"bff0000000");
KVEC(x"2",x"c0f0000000", x"40d0000000", x"bfd9999999");
KVEC(x"2",x"c0f0000000", x"40e0000000", x"bfcaaaaaaa");
KVEC(x"2",x"c0f0000000", x"40f0000000", x"bfc0000000");
KVEC(x"2",x"c0f0000000", x"4140000000", x"bf70000000");
KVEC(x"2",x"c0f0000000", x"4148000000", x"bf638e38e3");
KVEC(x"2",x"c0e0000000", x"c150000000", x"3f4ccccccc");
KVEC(x"2",x"c0e0000000", x"c148000000", x"3f55555555");
KVEC(x"2",x"c0e0000000", x"c140000000", x"3f60000000");
KVEC(x"5",x"0000000000", x"7fffffffff", x"7fffffffff");
KVEC(x"2",x"c0e0000000", x"c0f0000000", x"3f6db6db6c");
KVEC(x"2",x"c0e0000000", x"c0e0000000", x"3fc0000000");
KVEC(x"2",x"c0e0000000", x"c0d0000000", x"3fcccccccc");
KVEC(x"2",x"c0e0000000", x"c0c0000000", x"3fe0000000");
KVEC(x"2",x"c0e0000000", x"c060000000", x"4040000000");
KVEC(x"2",x"c0e0000000", x"c040000000", x"4060000000");
KVEC(x"2",x"c0e0000000", x"bfc0000000", x"40e0000000");
KVEC(x"2",x"c0e0000000", x"0000000000", x"ff80000000");
KVEC(x"2",x"c0e0000000", x"3fc0000000", x"c0e0000000");
KVEC(x"2",x"c0e0000000", x"4040000000", x"c060000000");
KVEC(x"5",x"7f80000000", x"40d0000000", x"7f80000000");
KVEC(x"2",x"c0e0000000", x"4060000000", x"c040000000");
KVEC(x"2",x"c0e0000000", x"40c0000000", x"bfe0000000");
KVEC(x"2",x"c0e0000000", x"40d0000000", x"bfcccccccc");
KVEC(x"2",x"c0e0000000", x"40e0000000", x"bfc0000000");
KVEC(x"2",x"c0e0000000", x"40f0000000", x"bf6db6db6c");
KVEC(x"2",x"c0e0000000", x"4140000000", x"bf60000000");
KVEC(x"2",x"c0e0000000", x"4148000000", x"bf55555555");
KVEC(x"2",x"c0d0000000", x"c150000000", x"3f40000000");
KVEC(x"2",x"c0d0000000", x"c148000000", x"3f471c71c7");
KVEC(x"2",x"c0d0000000", x"c140000000", x"3f50000000");
KVEC(x"5",x"7f80000000", x"0000000000", x"7f80000000");
KVEC(x"2",x"c0d0000000", x"c0f0000000", x"3f5b6db6da");
KVEC(x"2",x"c0d0000000", x"c0e0000000", x"3f6aaaaaaa");
KVEC(x"2",x"c0d0000000", x"c0d0000000", x"3fc0000000");
KVEC(x"2",x"c0d0000000", x"c0c0000000", x"3fd0000000");
KVEC(x"2",x"c0d0000000", x"c060000000", x"3feaaaaaaa");
KVEC(x"2",x"c0d0000000", x"c040000000", x"4050000000");
KVEC(x"2",x"c0d0000000", x"bfc0000000", x"40d0000000");
KVEC(x"2",x"c0d0000000", x"0000000000", x"ff80000000");
KVEC(x"2",x"c0d0000000", x"3fc0000000", x"c0d0000000");
KVEC(x"2",x"c0d0000000", x"4040000000", x"c050000000");
KVEC(x"5",x"7f80000000", x"7f80000000", x"7fffffffff");
KVEC(x"2",x"c0d0000000", x"4060000000", x"bfeaaaaaaa");
KVEC(x"2",x"c0d0000000", x"40c0000000", x"bfd0000000");
KVEC(x"2",x"c0d0000000", x"40d0000000", x"bfc0000000");
KVEC(x"2",x"c0d0000000", x"40e0000000", x"bf6aaaaaaa");
KVEC(x"2",x"c0d0000000", x"40f0000000", x"bf5b6db6da");
KVEC(x"2",x"c0d0000000", x"4140000000", x"bf50000000");
KVEC(x"2",x"c0d0000000", x"4148000000", x"bf471c71c7");
KVEC(x"2",x"c0c0000000", x"c150000000", x"3ee6666666");
KVEC(x"2",x"c0c0000000", x"c148000000", x"3ef1c71c70");
KVEC(x"2",x"c0c0000000", x"c140000000", x"3f40000000");
KVEC(x"5",x"7f80000000", x"ff80000000", x"7f80000000");
KVEC(x"2",x"c0c0000000", x"c0f0000000", x"3f49249248");
KVEC(x"2",x"c0c0000000", x"c0e0000000", x"3f55555554");
KVEC(x"2",x"c0c0000000", x"c0d0000000", x"3f66666666");
KVEC(x"2",x"c0c0000000", x"c0c0000000", x"3fc0000000");
KVEC(x"2",x"c0c0000000", x"c060000000", x"3fd5555554");
KVEC(x"2",x"c0c0000000", x"c040000000", x"4040000000");
KVEC(x"2",x"c0c0000000", x"bfc0000000", x"40c0000000");
KVEC(x"2",x"c0c0000000", x"0000000000", x"ff80000000");
KVEC(x"2",x"c0c0000000", x"3fc0000000", x"c0c0000000");
KVEC(x"2",x"c0c0000000", x"4040000000", x"c040000000");
KVEC(x"4",x"40d0000000", x"ff80000000", x"ff80000000");
KVEC(x"5",x"7f80000000", x"7fffffffff", x"7fffffffff");
KVEC(x"2",x"c0c0000000", x"4060000000", x"bfd5555554");
KVEC(x"2",x"c0c0000000", x"40c0000000", x"bfc0000000");
KVEC(x"2",x"c0c0000000", x"40d0000000", x"bf66666666");
KVEC(x"2",x"c0c0000000", x"40e0000000", x"bf55555554");
KVEC(x"2",x"c0c0000000", x"40f0000000", x"bf49249248");
KVEC(x"2",x"c0c0000000", x"4140000000", x"bf40000000");
KVEC(x"2",x"c0c0000000", x"4148000000", x"bef1c71c70");
KVEC(x"2",x"c060000000", x"c150000000", x"3ecccccccc");
KVEC(x"2",x"c060000000", x"c148000000", x"3ed5555555");
KVEC(x"2",x"c060000000", x"c140000000", x"3ee0000000");
KVEC(x"5",x"ff80000000", x"40d0000000", x"ff80000000");
KVEC(x"2",x"c060000000", x"c0f0000000", x"3eedb6db6c");
KVEC(x"2",x"c060000000", x"c0e0000000", x"3f40000000");
KVEC(x"2",x"c060000000", x"c0d0000000", x"3f4ccccccc");
KVEC(x"2",x"c060000000", x"c0c0000000", x"3f60000000");
KVEC(x"2",x"c060000000", x"c060000000", x"3fc0000000");
KVEC(x"2",x"c060000000", x"c040000000", x"3fe0000000");
KVEC(x"2",x"c060000000", x"bfc0000000", x"4060000000");
KVEC(x"2",x"c060000000", x"0000000000", x"ff80000000");
KVEC(x"2",x"c060000000", x"3fc0000000", x"c060000000");
KVEC(x"2",x"c060000000", x"4040000000", x"bfe0000000");
KVEC(x"5",x"ff80000000", x"0000000000", x"ff80000000");
KVEC(x"2",x"c060000000", x"4060000000", x"bfc0000000");
KVEC(x"2",x"c060000000", x"40c0000000", x"bf60000000");
KVEC(x"2",x"c060000000", x"40d0000000", x"bf4ccccccc");
KVEC(x"2",x"c060000000", x"40e0000000", x"bf40000000");
KVEC(x"2",x"c060000000", x"40f0000000", x"beedb6db6c");
KVEC(x"2",x"c060000000", x"4140000000", x"bee0000000");
KVEC(x"2",x"c060000000", x"4148000000", x"bed5555555");
KVEC(x"2",x"c040000000", x"c150000000", x"3e66666666");
KVEC(x"2",x"c040000000", x"c148000000", x"3e71c71c70");
KVEC(x"2",x"c040000000", x"c140000000", x"3ec0000000");
KVEC(x"5",x"ff80000000", x"7f80000000", x"ff80000000");
KVEC(x"2",x"c040000000", x"c0f0000000", x"3ec9249248");
KVEC(x"2",x"c040000000", x"c0e0000000", x"3ed5555554");
KVEC(x"2",x"c040000000", x"c0d0000000", x"3ee6666666");
KVEC(x"2",x"c040000000", x"c0c0000000", x"3f40000000");
KVEC(x"2",x"c040000000", x"c060000000", x"3f55555554");
KVEC(x"2",x"c040000000", x"c040000000", x"3fc0000000");
KVEC(x"2",x"c040000000", x"bfc0000000", x"4040000000");
KVEC(x"2",x"c040000000", x"0000000000", x"ff80000000");
KVEC(x"2",x"c040000000", x"3fc0000000", x"c040000000");
KVEC(x"2",x"c040000000", x"4040000000", x"bfc0000000");
KVEC(x"5",x"ff80000000", x"ff80000000", x"7fffffffff");
KVEC(x"2",x"c040000000", x"4060000000", x"bf55555554");
KVEC(x"2",x"c040000000", x"40c0000000", x"bf40000000");
KVEC(x"2",x"c040000000", x"40d0000000", x"bee6666666");
KVEC(x"2",x"c040000000", x"40e0000000", x"bed5555554");
KVEC(x"2",x"c040000000", x"40f0000000", x"bec9249248");
KVEC(x"2",x"c040000000", x"4140000000", x"bec0000000");
KVEC(x"2",x"c040000000", x"4148000000", x"be71c71c70");
KVEC(x"2",x"bfc0000000", x"c150000000", x"3de6666666");
KVEC(x"2",x"bfc0000000", x"c148000000", x"3df1c71c70");
KVEC(x"2",x"bfc0000000", x"c140000000", x"3e40000000");
KVEC(x"5",x"ff80000000", x"7fffffffff", x"7fffffffff");
KVEC(x"2",x"bfc0000000", x"c0f0000000", x"3e49249248");
KVEC(x"2",x"bfc0000000", x"c0e0000000", x"3e55555554");
KVEC(x"2",x"bfc0000000", x"c0d0000000", x"3e66666666");
KVEC(x"2",x"bfc0000000", x"c0c0000000", x"3ec0000000");
KVEC(x"2",x"bfc0000000", x"c060000000", x"3ed5555554");
KVEC(x"2",x"bfc0000000", x"c040000000", x"3f40000000");
KVEC(x"2",x"bfc0000000", x"bfc0000000", x"3fc0000000");
KVEC(x"2",x"bfc0000000", x"0000000000", x"ff80000000");
KVEC(x"2",x"bfc0000000", x"3fc0000000", x"bfc0000000");
KVEC(x"2",x"bfc0000000", x"4040000000", x"bf40000000");
KVEC(x"5",x"7fffffffff", x"40d0000000", x"7fffffffff");
KVEC(x"2",x"bfc0000000", x"4060000000", x"bed5555554");
KVEC(x"2",x"bfc0000000", x"40c0000000", x"bec0000000");
KVEC(x"2",x"bfc0000000", x"40d0000000", x"be66666666");
KVEC(x"2",x"bfc0000000", x"40e0000000", x"be55555554");
KVEC(x"2",x"bfc0000000", x"40f0000000", x"be49249248");
KVEC(x"2",x"bfc0000000", x"4140000000", x"be40000000");
KVEC(x"2",x"bfc0000000", x"4148000000", x"bdf1c71c70");
KVEC(x"2",x"0000000000", x"c150000000", x"8000000000");
KVEC(x"2",x"0000000000", x"c148000000", x"8000000000");
KVEC(x"2",x"0000000000", x"c140000000", x"8000000000");
KVEC(x"5",x"7fffffffff", x"0000000000", x"7fffffffff");
KVEC(x"2",x"0000000000", x"c0f0000000", x"8000000000");
KVEC(x"2",x"0000000000", x"c0e0000000", x"8000000000");
KVEC(x"2",x"0000000000", x"c0d0000000", x"8000000000");
KVEC(x"2",x"0000000000", x"c0c0000000", x"8000000000");
KVEC(x"2",x"0000000000", x"c060000000", x"8000000000");
KVEC(x"2",x"0000000000", x"c040000000", x"8000000000");
KVEC(x"2",x"0000000000", x"bfc0000000", x"8000000000");
KVEC(x"2",x"0000000000", x"0000000000", x"7fffffffff");
KVEC(x"2",x"0000000000", x"3fc0000000", x"0000000000");
KVEC(x"2",x"0000000000", x"4040000000", x"0000000000");
KVEC(x"5",x"7fffffffff", x"7f80000000", x"7fffffffff");
KVEC(x"2",x"0000000000", x"4060000000", x"0000000000");
KVEC(x"2",x"0000000000", x"40c0000000", x"0000000000");
KVEC(x"2",x"0000000000", x"40d0000000", x"0000000000");
KVEC(x"2",x"0000000000", x"40e0000000", x"0000000000");
KVEC(x"2",x"0000000000", x"40f0000000", x"0000000000");
KVEC(x"2",x"0000000000", x"4140000000", x"0000000000");
KVEC(x"2",x"0000000000", x"4148000000", x"0000000000");
KVEC(x"2",x"3fc0000000", x"c150000000", x"bde6666666");
KVEC(x"2",x"3fc0000000", x"c148000000", x"bdf1c71c70");
KVEC(x"2",x"3fc0000000", x"c140000000", x"be40000000");
KVEC(x"5",x"7fffffffff", x"ff80000000", x"7fffffffff");
KVEC(x"2",x"3fc0000000", x"c0f0000000", x"be49249248");
KVEC(x"2",x"3fc0000000", x"c0e0000000", x"be55555554");
KVEC(x"2",x"3fc0000000", x"c0d0000000", x"be66666666");
KVEC(x"2",x"3fc0000000", x"c0c0000000", x"bec0000000");
KVEC(x"2",x"3fc0000000", x"c060000000", x"bed5555554");
KVEC(x"2",x"3fc0000000", x"c040000000", x"bf40000000");
KVEC(x"2",x"3fc0000000", x"bfc0000000", x"bfc0000000");
KVEC(x"2",x"3fc0000000", x"0000000000", x"7f80000000");
KVEC(x"2",x"3fc0000000", x"3fc0000000", x"3fc0000000");
KVEC(x"2",x"3fc0000000", x"4040000000", x"3f40000000");
KVEC(x"4",x"40d0000000", x"7fffffffff", x"7fffffffff");
KVEC(x"5",x"7fffffffff", x"7fffffffff", x"7fffffffff");
KVEC(x"2",x"3fc0000000", x"4060000000", x"3ed5555554");
KVEC(x"2",x"3fc0000000", x"40c0000000", x"3ec0000000");
KVEC(x"2",x"3fc0000000", x"40d0000000", x"3e66666666");
KVEC(x"2",x"3fc0000000", x"40e0000000", x"3e55555554");
KVEC(x"2",x"3fc0000000", x"40f0000000", x"3e49249248");
KVEC(x"2",x"3fc0000000", x"4140000000", x"3e40000000");
KVEC(x"2",x"3fc0000000", x"4148000000", x"3df1c71c70");
KVEC(x"2",x"4040000000", x"c150000000", x"be66666666");
KVEC(x"2",x"4040000000", x"c148000000", x"be71c71c70");
KVEC(x"2",x"4040000000", x"c140000000", x"bec0000000");
KVEC(x"3",x"40d0000000", x"40d0000000", x"41e4000000");
KVEC(x"2",x"4040000000", x"c0f0000000", x"bec9249248");
KVEC(x"2",x"4040000000", x"c0e0000000", x"bed5555554");
KVEC(x"2",x"4040000000", x"c0d0000000", x"bee6666666");
KVEC(x"2",x"4040000000", x"c0c0000000", x"bf40000000");
KVEC(x"2",x"4040000000", x"c060000000", x"bf55555554");
KVEC(x"2",x"4040000000", x"c040000000", x"bfc0000000");
KVEC(x"2",x"4040000000", x"bfc0000000", x"c040000000");
KVEC(x"2",x"4040000000", x"0000000000", x"7f80000000");
KVEC(x"2",x"4040000000", x"3fc0000000", x"4040000000");
KVEC(x"2",x"4040000000", x"4040000000", x"3fc0000000");
KVEC(x"3",x"40d0000000", x"0000000000", x"0000000000");
KVEC(x"2",x"4040000000", x"4060000000", x"3f55555554");
KVEC(x"2",x"4040000000", x"40c0000000", x"3f40000000");
KVEC(x"2",x"4040000000", x"40d0000000", x"3ee6666666");
KVEC(x"2",x"4040000000", x"40e0000000", x"3ed5555554");
KVEC(x"2",x"4040000000", x"40f0000000", x"3ec9249248");
KVEC(x"2",x"4040000000", x"4140000000", x"3ec0000000");
KVEC(x"2",x"4040000000", x"4148000000", x"3e71c71c70");
KVEC(x"2",x"4060000000", x"c150000000", x"becccccccc");
KVEC(x"2",x"4060000000", x"c148000000", x"bed5555555");
KVEC(x"2",x"4060000000", x"c140000000", x"bee0000000");
KVEC(x"3",x"40d0000000", x"7f80000000", x"7f80000000");
KVEC(x"2",x"4060000000", x"c0f0000000", x"beedb6db6c");
KVEC(x"2",x"4060000000", x"c0e0000000", x"bf40000000");
KVEC(x"2",x"4060000000", x"c0d0000000", x"bf4ccccccc");
KVEC(x"2",x"4060000000", x"c0c0000000", x"bf60000000");
KVEC(x"2",x"4060000000", x"c060000000", x"bfc0000000");
KVEC(x"2",x"4060000000", x"c040000000", x"bfe0000000");
KVEC(x"2",x"4060000000", x"bfc0000000", x"c060000000");
KVEC(x"2",x"4060000000", x"0000000000", x"7f80000000");
KVEC(x"2",x"4060000000", x"3fc0000000", x"4060000000");
KVEC(x"2",x"4060000000", x"4040000000", x"3fe0000000");
KVEC(x"3",x"40d0000000", x"ff80000000", x"ff80000000");
KVEC(x"2",x"4060000000", x"4060000000", x"3fc0000000");
KVEC(x"2",x"4060000000", x"40c0000000", x"3f60000000");
KVEC(x"2",x"4060000000", x"40d0000000", x"3f4ccccccc");
KVEC(x"2",x"4060000000", x"40e0000000", x"3f40000000");
KVEC(x"2",x"4060000000", x"40f0000000", x"3eedb6db6c");
KVEC(x"2",x"4060000000", x"4140000000", x"3ee0000000");
KVEC(x"2",x"4060000000", x"4148000000", x"3ed5555555");
KVEC(x"2",x"40c0000000", x"c150000000", x"bee6666666");
KVEC(x"2",x"40c0000000", x"c148000000", x"bef1c71c70");
KVEC(x"2",x"40c0000000", x"c140000000", x"bf40000000");
KVEC(x"3",x"40d0000000", x"7fffffffff", x"7fffffffff");
KVEC(x"2",x"40c0000000", x"c0f0000000", x"bf49249248");
KVEC(x"2",x"40c0000000", x"c0e0000000", x"bf55555554");
KVEC(x"2",x"40c0000000", x"c0d0000000", x"bf66666666");
KVEC(x"2",x"40c0000000", x"c0c0000000", x"bfc0000000");
KVEC(x"2",x"40c0000000", x"c060000000", x"bfd5555554");
KVEC(x"2",x"40c0000000", x"c040000000", x"c040000000");
KVEC(x"2",x"40c0000000", x"bfc0000000", x"c0c0000000");
KVEC(x"2",x"40c0000000", x"0000000000", x"7f80000000");
KVEC(x"2",x"40c0000000", x"3fc0000000", x"40c0000000");
KVEC(x"2",x"40c0000000", x"4040000000", x"4040000000");
KVEC(x"3",x"0000000000", x"40d0000000", x"0000000000");
KVEC(x"2",x"40c0000000", x"4060000000", x"3fd5555554");
KVEC(x"2",x"40c0000000", x"40c0000000", x"3fc0000000");
KVEC(x"2",x"40c0000000", x"40d0000000", x"3f66666666");
KVEC(x"2",x"40c0000000", x"40e0000000", x"3f55555554");
KVEC(x"2",x"40c0000000", x"40f0000000", x"3f49249248");
KVEC(x"2",x"40c0000000", x"4140000000", x"3f40000000");
KVEC(x"2",x"40c0000000", x"4148000000", x"3ef1c71c70");
KVEC(x"2",x"40d0000000", x"c150000000", x"bf40000000");
KVEC(x"2",x"40d0000000", x"c148000000", x"bf471c71c7");
KVEC(x"2",x"40d0000000", x"c140000000", x"bf50000000");
KVEC(x"3",x"0000000000", x"0000000000", x"0000000000");
KVEC(x"2",x"40d0000000", x"c0f0000000", x"bf5b6db6da");
KVEC(x"2",x"40d0000000", x"c0e0000000", x"bf6aaaaaaa");
KVEC(x"2",x"40d0000000", x"c0d0000000", x"bfc0000000");
KVEC(x"2",x"40d0000000", x"c0c0000000", x"bfd0000000");
KVEC(x"2",x"40d0000000", x"c060000000", x"bfeaaaaaaa");
KVEC(x"2",x"40d0000000", x"c040000000", x"c050000000");
KVEC(x"2",x"40d0000000", x"bfc0000000", x"c0d0000000");
KVEC(x"2",x"40d0000000", x"0000000000", x"7f80000000");
KVEC(x"2",x"40d0000000", x"3fc0000000", x"40d0000000");
KVEC(x"2",x"40d0000000", x"4040000000", x"4050000000");
KVEC(x"3",x"0000000000", x"7f80000000", x"7fffffffff");
KVEC(x"2",x"40d0000000", x"4060000000", x"3feaaaaaaa");
KVEC(x"2",x"40d0000000", x"40c0000000", x"3fd0000000");
KVEC(x"2",x"40d0000000", x"40d0000000", x"3fc0000000");
KVEC(x"2",x"40d0000000", x"40e0000000", x"3f6aaaaaaa");
KVEC(x"2",x"40d0000000", x"40f0000000", x"3f5b6db6da");
KVEC(x"2",x"40d0000000", x"4140000000", x"3f50000000");
KVEC(x"2",x"40d0000000", x"4148000000", x"3f471c71c7");
KVEC(x"2",x"40e0000000", x"c150000000", x"bf4ccccccc");
KVEC(x"2",x"40e0000000", x"c148000000", x"bf55555555");
KVEC(x"2",x"40e0000000", x"c140000000", x"bf60000000");
KVEC(x"3",x"0000000000", x"ff80000000", x"7fffffffff");
KVEC(x"2",x"40e0000000", x"c0f0000000", x"bf6db6db6c");
KVEC(x"2",x"40e0000000", x"c0e0000000", x"bfc0000000");
KVEC(x"2",x"40e0000000", x"c0d0000000", x"bfcccccccc");
KVEC(x"2",x"40e0000000", x"c0c0000000", x"bfe0000000");
KVEC(x"2",x"40e0000000", x"c060000000", x"c040000000");
KVEC(x"2",x"40e0000000", x"c040000000", x"c060000000");
KVEC(x"2",x"40e0000000", x"bfc0000000", x"c0e0000000");
KVEC(x"2",x"40e0000000", x"0000000000", x"7f80000000");
KVEC(x"2",x"40e0000000", x"3fc0000000", x"40e0000000");
KVEC(x"2",x"40e0000000", x"4040000000", x"4060000000");
KVEC(x"4",x"0000000000", x"40d0000000", x"40d0000000");
KVEC(x"3",x"0000000000", x"7fffffffff", x"7fffffffff");
KVEC(x"2",x"40e0000000", x"4060000000", x"4040000000");
KVEC(x"2",x"40e0000000", x"40c0000000", x"3fe0000000");
KVEC(x"2",x"40e0000000", x"40d0000000", x"3fcccccccc");
KVEC(x"2",x"40e0000000", x"40e0000000", x"3fc0000000");
KVEC(x"2",x"40e0000000", x"40f0000000", x"3f6db6db6c");
KVEC(x"2",x"40e0000000", x"4140000000", x"3f60000000");
KVEC(x"2",x"40e0000000", x"4148000000", x"3f55555555");
KVEC(x"2",x"40f0000000", x"c150000000", x"bf59999999");
KVEC(x"2",x"40f0000000", x"c148000000", x"bf638e38e3");
KVEC(x"2",x"40f0000000", x"c140000000", x"bf70000000");
KVEC(x"3",x"7f80000000", x"40d0000000", x"7f80000000");
KVEC(x"2",x"40f0000000", x"c0f0000000", x"bfc0000000");
KVEC(x"2",x"40f0000000", x"c0e0000000", x"bfcaaaaaaa");
KVEC(x"2",x"40f0000000", x"c0d0000000", x"bfd9999999");
KVEC(x"2",x"40f0000000", x"c0c0000000", x"bff0000000");
KVEC(x"2",x"40f0000000", x"c060000000", x"c04aaaaaaa");
KVEC(x"2",x"40f0000000", x"c040000000", x"c070000000");
KVEC(x"2",x"40f0000000", x"bfc0000000", x"c0f0000000");
KVEC(x"2",x"40f0000000", x"0000000000", x"7f80000000");
KVEC(x"2",x"40f0000000", x"3fc0000000", x"40f0000000");
KVEC(x"2",x"40f0000000", x"4040000000", x"4070000000");
KVEC(x"3",x"7f80000000", x"0000000000", x"7fffffffff");
KVEC(x"2",x"40f0000000", x"4060000000", x"404aaaaaaa");
KVEC(x"2",x"40f0000000", x"40c0000000", x"3ff0000000");
KVEC(x"2",x"40f0000000", x"40d0000000", x"3fd9999999");
KVEC(x"2",x"40f0000000", x"40e0000000", x"3fcaaaaaaa");
KVEC(x"2",x"40f0000000", x"40f0000000", x"3fc0000000");
KVEC(x"2",x"40f0000000", x"4140000000", x"3f70000000");
KVEC(x"2",x"40f0000000", x"4148000000", x"3f638e38e3");
KVEC(x"2",x"4140000000", x"c150000000", x"bf66666666");
KVEC(x"2",x"4140000000", x"c148000000", x"bf71c71c70");
KVEC(x"2",x"4140000000", x"c140000000", x"bfc0000000");
KVEC(x"3",x"7f80000000", x"7f80000000", x"7f80000000");
KVEC(x"2",x"4140000000", x"c0f0000000", x"bfc9249248");
KVEC(x"2",x"4140000000", x"c0e0000000", x"bfd5555554");
KVEC(x"2",x"4140000000", x"c0d0000000", x"bfe6666666");
KVEC(x"2",x"4140000000", x"c0c0000000", x"c040000000");
KVEC(x"2",x"4140000000", x"c060000000", x"c055555554");
KVEC(x"2",x"4140000000", x"c040000000", x"c0c0000000");
KVEC(x"2",x"4140000000", x"bfc0000000", x"c140000000");
KVEC(x"2",x"4140000000", x"0000000000", x"7f80000000");
KVEC(x"2",x"4140000000", x"3fc0000000", x"4140000000");
KVEC(x"2",x"4140000000", x"4040000000", x"40c0000000");
KVEC(x"3",x"7f80000000", x"ff80000000", x"ff80000000");
KVEC(x"2",x"4140000000", x"4060000000", x"4055555554");
KVEC(x"2",x"4140000000", x"40c0000000", x"4040000000");
KVEC(x"2",x"4140000000", x"40d0000000", x"3fe6666666");
KVEC(x"2",x"4140000000", x"40e0000000", x"3fd5555554");
KVEC(x"2",x"4140000000", x"40f0000000", x"3fc9249248");
KVEC(x"2",x"4140000000", x"4140000000", x"3fc0000000");
KVEC(x"2",x"4140000000", x"4148000000", x"3f71c71c70");
KVEC(x"2",x"4148000000", x"c150000000", x"bf73333332");
KVEC(x"2",x"4148000000", x"c148000000", x"bfc0000000");
KVEC(x"2",x"4148000000", x"c140000000", x"bfc8000000");
KVEC(x"3",x"7f80000000", x"7fffffffff", x"7fffffffff");
KVEC(x"2",x"4148000000", x"c0f0000000", x"bfd2492492");
KVEC(x"2",x"4148000000", x"c0e0000000", x"bfe0000000");
KVEC(x"2",x"4148000000", x"c0d0000000", x"bff3333332");
KVEC(x"2",x"4148000000", x"c0c0000000", x"c048000000");
KVEC(x"2",x"4148000000", x"c060000000", x"c060000000");
KVEC(x"2",x"4148000000", x"c040000000", x"c0c8000000");
KVEC(x"2",x"4148000000", x"bfc0000000", x"c148000000");
KVEC(x"2",x"4148000000", x"0000000000", x"7f80000000");
KVEC(x"2",x"4148000000", x"3fc0000000", x"4148000000");
KVEC(x"2",x"4148000000", x"4040000000", x"40c8000000");
KVEC(x"3",x"ff80000000", x"40d0000000", x"ff80000000");
KVEC(x"2",x"4148000000", x"4060000000", x"4060000000");
KVEC(x"2",x"4148000000", x"40c0000000", x"4048000000");
KVEC(x"2",x"4148000000", x"40d0000000", x"3ff3333332");
KVEC(x"2",x"4148000000", x"40e0000000", x"3fe0000000");
KVEC(x"2",x"4148000000", x"40f0000000", x"3fd2492492");
KVEC(x"2",x"4148000000", x"4140000000", x"3fc8000000");
KVEC(x"2",x"4148000000", x"4148000000", x"3fc0000000");
KVEC(x"3",x"0000000000", x"4178000000", x"0000000000");
KVEC(x"3",x"4178000000", x"0000000000", x"0000000000");
KVEC(x"3",x"4178000000", x"3fc0000000", x"4178000000");
KVEC(x"3",x"ff80000000", x"0000000000", x"7fffffffff");
KVEC(x"3",x"c178000000", x"4168000000", x"c361800000");
KVEC(x"3",x"4178000000", x"c168000000", x"c361800000");
KVEC(x"3",x"ce77359400", x"4e79a13564", x"dd7146c905");
KVEC(x"3",x"4178000000", x"7fffffffff", x"7fffffffff");
KVEC(x"3",x"7fffffffff", x"4178000000", x"7fffffffff");
KVEC(x"3",x"7fffffffff", x"7fffffffff", x"7fffffffff");
KVEC(x"4",x"0000000000", x"0000000000", x"0000000000");
KVEC(x"4",x"40e0000000", x"0000000000", x"40e0000000");
KVEC(x"4",x"0000000000", x"40e0000000", x"40e0000000");
KVEC(x"4",x"40d0000000", x"40c0000000", x"4148000000");
KVEC(x"3",x"ff80000000", x"7f80000000", x"ff80000000");
KVEC(x"4",x"40d0000000", x"c0c0000000", x"3fc0000000");
KVEC(x"4",x"c0d0000000", x"40c0000000", x"bfc0000000");
KVEC(x"4",x"c0d0000000", x"c0c0000000", x"c148000000");
KVEC(x"5",x"35c31bde82", x"33eb5fca6a", x"3578cbc3b8");
KVEC(x"5",x"35c31bde82", x"12cf3a68db", x"35c31bde82");
KVEC(x"5",x"0000000000", x"0000000000", x"0000000000");
KVEC(x"5",x"40e0000000", x"0000000000", x"40e0000000");
KVEC(x"5",x"0000000000", x"40e0000000", x"c0e0000000");
KVEC(x"5",x"4148000000", x"40c0000000", x"40d0000000");
KVEC(x"5",x"4148000000", x"c0c0000000", x"4168000000");
KVEC(x"3",x"ff80000000", x"ff80000000", x"7f80000000");
KVEC(x"5",x"c148000000", x"40c0000000", x"c168000000");
KVEC(x"5",x"c148000000", x"c0c0000000", x"c0d0000000");
KVEC(x"5",x"35c31bde82", x"33eb5fca6a", x"3578cbc3b8");
KVEC(x"5",x"35c31bde82", x"12cf3a68db", x"35c31bde82");
KVEC(x"4",x"0000000000", x"0000000000", x"0000000000");
KVEC(x"3",x"ff80000000", x"7fffffffff", x"7fffffffff");
KVEC(x"3",x"7fffffffff", x"40d0000000", x"7fffffffff");
KVEC(x"3",x"7fffffffff", x"0000000000", x"7fffffffff");
KVEC(x"3",x"7fffffffff", x"7f80000000", x"7fffffffff");
KVEC(x"3",x"7fffffffff", x"ff80000000", x"7fffffffff");
KVEC(x"3",x"7fffffffff", x"7fffffffff", x"7fffffffff");
KVEC(x"2",x"40d0000000", x"40d0000000", x"3fc0000000");
KVEC(x"2",x"40d0000000", x"0000000000", x"7f80000000");
KVEC(x"2",x"40d0000000", x"7f80000000", x"0000000000");
KVEC(x"2",x"40d0000000", x"ff80000000", x"8000000000");
KVEC(x"4",x"0000000000", x"7f80000000", x"7f80000000");
KVEC(x"2",x"40d0000000", x"7fffffffff", x"7fffffffff");
KVEC(x"2",x"0000000000", x"40d0000000", x"0000000000");
KVEC(x"2",x"0000000000", x"0000000000", x"7fffffffff");
KVEC(x"2",x"0000000000", x"7f80000000", x"0000000000");
KVEC(x"2",x"0000000000", x"ff80000000", x"8000000000");
KVEC(x"2",x"0000000000", x"7fffffffff", x"7fffffffff");
KVEC(x"2",x"7f80000000", x"40d0000000", x"7f80000000");
KVEC(x"2",x"7f80000000", x"0000000000", x"7f80000000");
KVEC(x"2",x"7f80000000", x"7f80000000", x"7fffffffff");
KVEC(x"2",x"7f80000000", x"ff80000000", x"7fffffffff");
KVEC(x"4",x"0000000000", x"ff80000000", x"ff80000000");
KVEC(x"2",x"7f80000000", x"7fffffffff", x"7fffffffff");
KVEC(x"2",x"ff80000000", x"40d0000000", x"ff80000000");
KVEC(x"2",x"ff80000000", x"0000000000", x"ff80000000");
KVEC(x"2",x"ff80000000", x"7f80000000", x"7fffffffff");
KVEC(x"2",x"ff80000000", x"ff80000000", x"7fffffffff");
KVEC(x"2",x"ff80000000", x"7fffffffff", x"7fffffffff");
KVEC(x"2",x"7fffffffff", x"40d0000000", x"7fffffffff");
KVEC(x"2",x"7fffffffff", x"0000000000", x"7fffffffff");
KVEC(x"2",x"7fffffffff", x"7f80000000", x"7fffffffff");
KVEC(x"2",x"7fffffffff", x"ff80000000", x"7fffffffff");

    err_count := 0;


    -- we have 8 bits of precision in the output, so if we use
    -- really large periods we're going to lose significant figures
    -- and be totally inaccurate, so we only go close to top end
    per := 100;
    while per < 2 ** (32-8) loop
      run_uint( "0000", 1000000000, per);
      per := per + 100 + per/10;
    end loop;



    simulation_done <= true;

    report "KMATH Complete: " & integer'image(failures) & " failures, " &
      integer'image(err_count) & " out of range warnings, " &
      integer'image(vec_fails) & " vector fails " &
      " in " &
      integer'image(runs) & " runs.";

    wait;                               -- till the end of time

  end process p;


end Behavioral;
